`timescale 1ns/1ns

`include "../src/riscv_core/opcode.vh"
`include "mem_path.vh"

// This testbench tests if the cpu module can decode and execute
// all the instructions specified in the spec (RV32I -- including CSRRW and CSRRWI).
// Some tests for data hazards and control hazards are also included.

// How does the testbench work?
// For each test, the testbench initializes IMem with one or several instructions
// (encoded in binary format as specified in the spec) for testing.
// RegFile and DMem are also initialized with some data.
// Then, the clock is advanced until the cpu module gives correct result
// in the RegFile or DMem. If no correct result is returned after a "timeout" cycle,
// the testbench will be terminated (or failed)

// This setting is different from other testbenches, in which the BIOSMem or IMem is initialized
// with a hex file generated by compiling the assembly/C code of the corresponding
// test software (the hex file contains the binary encoding of the instructions and data
// of the program). Here, we manually generate the instructions and data.

// Don't just run the testbench, look at the tests, see what they do.
// The testbench is intended to provide you some examples to get started.
// Feel free to make your own change.
// Note that the testbench is by no means exhaustive.
// You should add your own tests if there are cases you think the testbench
// does not cover.

module fpu_tb();
  reg clk, rst;
  parameter CPU_CLOCK_PERIOD = 20;
  parameter CPU_CLOCK_FREQ   = 1_000_000_000 / CPU_CLOCK_PERIOD;

  initial clk = 0;
  always #(CPU_CLOCK_PERIOD/2) clk = ~clk;
  wire [31:0] csr;
  reg bp_enable = 1'b0;

  // Init PC with 32'h1000_0000 -- address space of IMem
  // When PC is in IMem's address space, IMem is read-only
  // DMem can be R/W as long as the addr bits [31:28] is 4'b00x1
  cpu # (
    .CPU_CLOCK_FREQ(CPU_CLOCK_FREQ),
    .RESET_PC(32'h1000_0000)
  ) cpu (
    .clk(clk),
    .rst(rst),
    .bp_enable(bp_enable),
    .serial_in(1'b1),
    .serial_out()
  );

  wire [31:0] timeout_cycle = 1000;

  // Reset IMem, DMem, and RegFile before running new test
  task reset;
    integer i;
    begin
      for (i = 0; i < `RF_PATH.DEPTH; i = i + 1) begin
        `RF_PATH.mem[i] = 0;
        `FPRF_PATH.mem[i] = 0;
      end
      for (i = 0; i < `DMEM_PATH.DEPTH; i = i + 1) begin
        `DMEM_PATH.mem[i] = 0;
      end
      for (i = 0; i < `IMEM_PATH.DEPTH; i = i + 1) begin
        `IMEM_PATH.mem[i] = 0;
      end
    end
  endtask

  task reset_cpu;
    @(negedge clk);
    rst = 1;
    @(negedge clk);
    rst = 0;
  endtask

  task init_rf;
    integer i;
    begin
      for (i = 1; i < `RF_PATH.DEPTH; i = i + 1) begin
        `RF_PATH.mem[i] = 100 * i + 1;
      end
    end
  endtask

  reg [31:0] cycle;
  reg done;
  reg [31:0]  current_test_id = 0;
  reg [255:0] current_test_type;
  reg [31:0]  current_output;
  reg [31:0]  current_result;
  reg all_tests_passed = 0;


  // Check for timeout
  // If a test does not return correct value in a given timeout cycle,
  // we terminate the testbench
  initial begin
    while (all_tests_passed === 0) begin
      @(posedge clk);
      if (cycle === timeout_cycle) begin
        $display("[Failed] Timeout at [%d] test %s, expected_result = %h, got = %h",
                current_test_id, current_test_type, current_result, current_output);
        $finish();
      end
    end
  end

  always @(posedge clk) begin
    if (done === 0)
      cycle <= cycle + 1;
    else
      cycle <= 0;
  end

  // Check result of RegFile
  // If the write_back (destination) register has correct value (matches "result"), test passed
  // This is used to test instructions that update RegFile
  task check_result_rf;
    input [31:0]  rf_wa;
    input [31:0]  result;
    input [255:0] test_type;
    begin
      done = 0;
      current_test_id   = current_test_id + 1;
      current_test_type = test_type;
      current_result    = result;
      while (`RF_PATH.mem[rf_wa] !== result) begin
        current_output = `RF_PATH.mem[rf_wa];
        @(posedge clk);
      end
      cycle = 0;
      done = 1;
      $display("[%d] Test %s passed!", current_test_id, test_type);
    end
  endtask

  task check_result_fprf;
    input [31:0]  rf_wa;
    input [31:0]  result;
    input [255:0] test_type;
    begin
      done = 0;
      current_test_id   = current_test_id + 1;
      current_test_type = test_type;
      current_result    = result;
      while (`FPRF_PATH.mem[rf_wa] !== result) begin
        current_output = `FPRF_PATH.mem[rf_wa];
        @(posedge clk);
      end
      cycle = 0;
      done = 1;
      $display("[%d] Test %s passed!", current_test_id, test_type);
    end
  endtask

  // Check result of DMem
  // If the memory location of DMem has correct value (matches "result"), test passed
  // This is used to test store instructions
  task check_result_dmem;
    input [31:0]  addr;
    input [31:0]  result;
    input [255:0] test_type;
    begin
      done = 0;
      current_test_id   = current_test_id + 1;
      current_test_type = test_type;
      current_result    = result;
      while (`DMEM_PATH.mem[addr] !== result) begin
        current_output = `DMEM_PATH.mem[addr];
        @(posedge clk);
      end
      cycle = 0;
      done = 1;
      $display("[%d] Test %s passed!", current_test_id, test_type);
    end
  endtask

  integer i;

  reg [31:0] num_cycles = 0;
  reg [31:0] num_insts  = 0;
  reg [4:0]  RD, RS1, RS2, RS3;
  reg [31:0] RD1, RD2, RD3;
  reg [4:0]  SHAMT;
  reg [31:0] IMM, IMM0, IMM1, IMM2, IMM3;
  reg [14:0] INST_ADDR;
  reg [14:0] DATA_ADDR;
  reg [14:0] DATA_ADDR0, DATA_ADDR1, DATA_ADDR2, DATA_ADDR3;
  reg [14:0] DATA_ADDR4, DATA_ADDR5, DATA_ADDR6, DATA_ADDR7;
  reg [14:0] DATA_ADDR8, DATA_ADDR9;

  reg [31:0] JUMP_ADDR;

  reg [31:0]  BR_TAKEN_OP1  [5:0];
  reg [31:0]  BR_TAKEN_OP2  [5:0];
  reg [31:0]  BR_NTAKEN_OP1 [5:0];
  reg [31:0]  BR_NTAKEN_OP2 [5:0];
  reg [2:0]   BR_TYPE       [5:0];
  reg [255:0] BR_NAME_TK1   [5:0];
  reg [255:0] BR_NAME_TK2   [5:0];
  reg [255:0] BR_NAME_NTK   [5:0];

  initial begin
    `ifndef IVERILOG
        $vcdpluson;
    `endif
    `ifdef IVERILOG
        $dumpfile("cpu_tb.fst");
        $dumpvars(0, cpu_tb);
    `endif

    #0;
    rst = 0;

    // Reset the CPU
    rst = 1;
    // Hold reset for a while
    repeat (10) @(posedge clk);

    @(negedge clk);
    rst = 0;

    reset();

    // We can also use $random to generate random values for testing
    RS1 = 1; RD1 = 32'h400ccccd;
    RS2 = 2; RD2 = 32'h400ccccd;
    RS3 = 3; RD3 = 32'hbf570a3d;
    `FPRF_PATH.mem[RS1] = RD1; // 2.2
    `FPRF_PATH.mem[RS2] = RD2; // 2.2
    `FPRF_PATH.mem[RS3] = RD3; // 2.2
    `FPRF_PATH.mem[5'd21] = 32'h410d70a4; // 8.84
    `FPRF_PATH.mem[5'd22] = 32'hbf570a3d; // -.84
    `FPRF_PATH.mem[5'd29] = 32'h408ccccd; // 4.4
    `FPRF_PATH.mem[5'd30] = 32'h400ccccd; // 2.2
    `FPRF_PATH.mem[5'd31] = 32'hbf570a3d; // -.84
    `FPRF_PATH.mem[5'd18] = 32'hBf800000; // -1
    `FPRF_PATH.mem[5'd19] = 32'h40000000; // 2

    `RF_PATH.mem[5'd15] = 32'hDEADBEEF;
    `RF_PATH.mem[5'd16] = 32'd15;
    `RF_PATH.mem[5]  = 32'h3150_4000;
    `RF_PATH.mem[7]  = 32'h3150_8000;
    SHAMT           = 5'd20;
    INST_ADDR       = 14'h0000;

    `IMEM_PATH.mem[INST_ADDR] = 32'h0020F253; // fadd.s f4 f1 f2
    `IMEM_PATH.mem[INST_ADDR + 1] = 32'h1820F2C3; // fmadd.s f5, f1, f2, f3
    `IMEM_PATH.mem[INST_ADDR + 2] = 32'he0008353; // fmv.x.w x6 f1
    `IMEM_PATH.mem[INST_ADDR + 3] = 32'hF00783D3; // fmv.w.x f7 x15
    `IMEM_PATH.mem[INST_ADDR + 4] = 32'hD0087453; // fcvt.s.w f8 x16
    `IMEM_PATH.mem[INST_ADDR + 5] = 32'h203104d3; // fsgnj.s f9 f2 f3
    `IMEM_PATH.mem[INST_ADDR + 6] = 32'h0002a507; // flw f10 0(x5)
    `IMEM_PATH.mem[INST_ADDR + 7] = 32'h00a3a027; // fsw f10 0(x7)
    `IMEM_PATH.mem[INST_ADDR + 8] = 32'h013978d3; // fadd.s f17 f18 f19
    `IMEM_PATH.mem[INST_ADDR + 9] = 32'h016afa53; // fadd.s f20 f21 f22
    `IMEM_PATH.mem[INST_ADDR + 10] = 32'hf9eefe43; // fmadd.s f28 f29 f30 f31

    `DMEM_PATH.mem[14'h1000] = 32'hDEADBEEF;
    `DMEM_PATH.mem[14'h2000] = 32'h0;

    reset_cpu();

    check_result_fprf(5'd4,  32'h408ccccd, "FADD");
    check_result_fprf(5'd5,  32'h40800000, "FMADD");
    check_result_rf(5'd6, 32'h400ccccd, "FMV.X.W");
    check_result_fprf(5'd7,  32'hDEADBEEF, "FMV.W.X");
    check_result_fprf(5'd8, 32'h41700000, "FCVT.S.W");
    check_result_fprf(5'd9, 32'hc00ccccd, "FSGNJ.S");
    check_result_fprf(32'd10, 32'hDEADBEEF, "FLW");
    check_result_dmem(14'h2000, 32'hDEADBEEF, "FSW");
    check_result_fprf(5'd17,  32'h3f800000, "FADD - 2");
    check_result_fprf(5'd20,  32'h41000000, "FADD - 3");
    check_result_fprf(5'd28,  32'h410d70a4, "FMADD - 2");

    reset();

    // We can also use $random to generate random values for testing
    RS1 = 1; RD1 = 32'h400ccccd;  // 2.2
    RS2 = 2; RD2 = 32'h400ccccd;  // 2.2
    RS3 = 3; RD3 = 32'hbf570a3d;  // -.84
    `FPRF_PATH.mem[RS1] = RD1;
    `FPRF_PATH.mem[RS2] = RD2;
    `FPRF_PATH.mem[RS3] = RD3;
    `FPRF_PATH.mem[5'd4]=0;
    `FPRF_PATH.mem[5'd5]=0;


    SHAMT           = 5'd20;
    INST_ADDR       = 14'h0000;

    `IMEM_PATH.mem[INST_ADDR]  = 32'h0020F253; // fadd.s f4 f1 f2 ((2.2 + 2.2) * 2.2) - .84 = (4.4 * 2.2) - .84 = 9.68 -.84 = 8.84
    `IMEM_PATH.mem[INST_ADDR + 1]  = 32'h182272c3; // fmadd.s f5, f4, f2, f3

    reset_cpu();

    check_result_fprf(5'd4,  32'h408ccccd, "FADD -> FMADD hazard - 1");
    check_result_fprf(5'd5,  32'h410d70a4, "FADD -> FMADD hazard - 2");

    reset();

    // We can also use $random to generate random values for testing
    RS1 = 1; RD1 = 32'h400ccccd;
    RS2 = 2; RD2 = 32'h400ccccd;
    RS3 = 3; RD3 = 32'hbf570a3d; // -2.2
    `FPRF_PATH.mem[RS1] = RD1;
    `FPRF_PATH.mem[RS2] = RD2;
    `FPRF_PATH.mem[RS3] = RD3;
    SHAMT           = 5'd20;
    INST_ADDR       = 14'h0000;

    `IMEM_PATH.mem[INST_ADDR]  = 32'h1820f2c3; // fmadd.s f5, f1, f2, f3
    `IMEM_PATH.mem[INST_ADDR + 1]  = 32'h0022F253; // fadd.s f4 f5 f2

    reset_cpu();

    check_result_fprf(5'd5,  32'h40800000, "FMADD -> FADD hazard - 1");
    check_result_fprf(5'd4,  32'h40c66666, "FMADD -> FADD hazard - 2");



    all_tests_passed = 1'b1;

    repeat (100) @(posedge clk);
    $display("All tests passed!");
    $finish();
  end

endmodule